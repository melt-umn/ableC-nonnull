grammar edu:umn:cs:melt:exts:ableC:nonnull:src ;

exports edu:umn:cs:melt:exts:ableC:nonnull:src:abstractsyntax ;
exports edu:umn:cs:melt:exts:ableC:nonnull:src:concretesyntax ;

