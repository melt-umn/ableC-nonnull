grammar edu:umn:cs:melt:exts:ableC:nonnull:src:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:nonnull:src:concretesyntax:typeQualifier;


