grammar edu:umn:cs:melt:exts:ableC:nonnull;

exports edu:umn:cs:melt:exts:ableC:nonnull:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:nonnull:concretesyntax;

