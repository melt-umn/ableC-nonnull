grammar edu:umn:cs:melt:exts:ableC:nonnull:modular_analyses:determinism;

import edu:umn:cs:melt:ableC:host only ablecParser;

copper_mda testTypeQualifier(ablecParser) {
  edu:umn:cs:melt:exts:ableC:nonnull:src:concretesyntax:typeQualifier;
}

